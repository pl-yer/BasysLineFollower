

 module PID_controller(
    
    );
endmodule